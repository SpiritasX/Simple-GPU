library ieee;
use ieee.std_logic_1164.all;

library work;

entity gpu is
	Port (
		
	);
end gpu;

architecture Behavioral of gpu
	
begin
	
end Behavioral;