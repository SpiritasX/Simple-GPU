library ieee;
use ieee.std_logic_1164.all;

entity gpu_top is
	Port (
		
	);
end gpu_top;

architecture Behavioral of gpu_top
begin
	
end Behavioral;